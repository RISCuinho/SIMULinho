module SIMULinho;
initial $hello;
endmodule
