module SIMULinho;
initial begin
#1 $hello;
#2 $openUI;
#500 $closeUI;
end

endmodule
